library ieee;
use ieee.std_logic_1164.all;

entity main is
end entity;

architecture sim of main is

begin


end process;



end architecture;
